----------------------------------------------------------------------------------
-- COMPANY:		Ruhr University Bochum, Embedded Security
-- AUTHOR:		https://eprint.iacr.org/2018/203
----------------------------------------------------------------------------------
-- Copyright (c) 2019, Amir Moradi, Aein Rezaei Shahmirzadi
-- All rights reserved.

-- BSD-3-Clause License
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--     * Redistributions of source code must retain the above copyright
--       notice, this list of conditions and the following disclaimer.
--     * Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
--     * Neither the name of the copyright holder, their organization nor the
--       names of its contributors may be used to endorse or promote products
--       derived from this software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY F8 IS
	GENERIC ( size  : POSITIVE := 8;
				 count : POSITIVE; 
	          Table : STD_LOGIC_VECTOR (4095 DOWNTO 0));
	PORT ( data_in:  IN  STD_LOGIC_VECTOR (size*count-1    DOWNTO 0);
			 data_out: OUT STD_LOGIC_VECTOR (size*count-1 DOWNTO 0));
END F8;

ARCHITECTURE behavioral OF F8 IS
		SIGNAL CompressedData : STD_LOGIC_VECTOR(8*count-1 DOWNTO 0);
BEGIN

	CompressData_Inst: ENTITY work.CompressData
	GENERIC Map ( Red_size => size, count => count)
	PORT MAP(
		x  => data_in,
		y => CompressedData);
		
	GEN :
	FOR i IN 0 TO count-1 GENERATE
		LookUpSizex256_Inst: ENTITY work.LookUpSizex256
		Generic Map ( size, Table)
		Port Map (
			input		=> CompressedData ((i+1)*8-1    downto i*8),
			output	=> data_out((i+1)*size-1 downto i*size)
			);
			
	END GENERATE;
			
END behavioral;



