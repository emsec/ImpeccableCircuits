----------------------------------------------------------------------------------
-- COMPANY:		Ruhr University Bochum, Embedded Security
-- AUTHOR:		https://eprint.iacr.org/2018/203
----------------------------------------------------------------------------------
-- Copyright (c) 2019, Anita Aghaie, Amir Moradi, Aein Rezaei Shahmirzadi
-- All rights reserved.

-- BSD-3-Clause License
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--     * Redistributions of source code must retain the above copyright
--       notice, this list of conditions and the following disclaimer.
--     * Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
--     * Neither the name of the copyright holder, their organization nor the
--       names of its contributors may be used to endorse or promote products
--       derived from this software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity RedFinalRoundControlLogic is
    Generic ( 
		Red_size			: NATURAL;
		LFTable    		: STD_LOGIC_VECTOR (4095 DOWNTO 0);
		LFInvTable    		: STD_LOGIC_VECTOR (4095 DOWNTO 0));
   Port ( 
		Red_rcon   					: in   STD_LOGIC_VECTOR (Red_size-1 downto 0);
		Red_FinalRoundBit		: out  STD_LOGIC_VECTOR (Red_size-1 downto 0));
end RedFinalRoundControlLogic;

architecture Behavioral of RedFinalRoundControlLogic is
begin

	GEN :
	FOR i IN 0 TO Red_size-1 GENERATE
	
		RedFinalRoundControlLogicBit_Inst: ENTITY work.RedFinalRoundControlLogicBit 
		Generic Map (Red_size, LFTable, LFInvTable, i)
		PORT MAP(
			Red_rcon 			=> Red_rcon,
			Red_FinalRoundBit => Red_FinalRoundBit(i));
			
	END GENERATE;

end Behavioral;

