----------------------------------------------------------------------------------
-- COMPANY:		Ruhr University Bochum, Embedded Security
-- AUTHOR:		https://eprint.iacr.org/2018/203
----------------------------------------------------------------------------------
-- Copyright (c) 2019, Anita Aghaie, Amir Moradi
-- All rights reserved.

-- BSD-3-Clause License
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--     * Redistributions of source code must retain the above copyright
--       notice, this list of conditions and the following disclaimer.
--     * Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
--     * Neither the name of the copyright holder, their organization nor the
--       names of its contributors may be used to endorse or promote products
--       derived from this software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.functions.all;

-- Red_size     : 1 => LF: 0110100110010110
-- Red_size     : 2 => LF: 0132231032011023
-- Red_size     : 3 => LF: 0374562165123047

-- MultiVariate : 0 => Univariate   adversary model
-- MultiVariate : 1 => Multivariate adversary model

entity LED128Enc is
	 Generic ( Red_size  : POSITIVE := 1;
		   LFC       : STD_LOGIC_VECTOR (3  DOWNTO 0) := x"0";
	           LF        : STD_LOGIC_VECTOR (63 DOWNTO 0) := x"0110100110010110";
		   MultiVariate : NATURAL  := 0);
    Port ( clk 			: in  STD_LOGIC;
           rst 			: in  STD_LOGIC;
           Plaintext 	: in  STD_LOGIC_VECTOR ( 63 downto 0);
           Key 			: in  STD_LOGIC_VECTOR (127 downto 0);
           Ciphertext 	: out STD_LOGIC_VECTOR ( 63 downto 0);
           done 			: out STD_LOGIC);
end LED128Enc;

architecture Behavioral of LED128Enc is

	constant SboxTable : STD_LOGIC_VECTOR (63 DOWNTO 0) := x"C56B90AD3EF84712";

	constant LFTable   : STD_LOGIC_VECTOR (63 DOWNTO 0) := 
		(LF(63 downto 60) XOR LFC) &
		(LF(59 downto 56) XOR LFC) &
		(LF(55 downto 52) XOR LFC) &
		(LF(51 downto 48) XOR LFC) &
		(LF(47 downto 44) XOR LFC) &
		(LF(43 downto 40) XOR LFC) &
		(LF(39 downto 36) XOR LFC) &
		(LF(35 downto 32) XOR LFC) &
		(LF(31 downto 28) XOR LFC) &
		(LF(27 downto 24) XOR LFC) &
		(LF(23 downto 20) XOR LFC) &
		(LF(19 downto 16) XOR LFC) &
		(LF(15 downto 12) XOR LFC) &
		(LF(11 downto  8) XOR LFC) &
		(LF( 7 downto  4) XOR LFC) &
		(LF( 3 downto  0) XOR LFC);
	
	constant Identity : STD_LOGIC_VECTOR (63 DOWNTO 0) := x"0123456789ABCDEF";
	
	constant ToCheckCount : NATURAL := 5+16+18*MultiVariate;

	constant Distance 	 : NATURAL := GetDistance(Red_size, LFTable);
	constant Error_size   : NATURAL := Distance-1+Distance*MultiVariate;
	
	-------------------------------

	signal StateRegInput 						: STD_LOGIC_VECTOR(63 downto 0);
	signal StateRegOutput						: STD_LOGIC_VECTOR(63 downto 0);
	signal AddRoundKeyOutput					: STD_LOGIC_VECTOR(63 downto 0);
	signal AddKeyMUXOutput						: STD_LOGIC_VECTOR(63 downto 0);
	signal AddConstInput							: STD_LOGIC_VECTOR(31 downto 0);
	signal AddConstInput2						: STD_LOGIC_VECTOR(7  downto 0);
	signal AddConstOutput						: STD_LOGIC_VECTOR(31 downto 0);
	signal AddconstMUXOutput					: STD_LOGIC_VECTOR(31 downto 0);
	signal ShiftRowsInput						: STD_LOGIC_VECTOR(63 downto 0);
	signal ShiftRowsOutput						: STD_LOGIC_VECTOR(63 downto 0);
	signal Feedback								: STD_LOGIC_VECTOR(63 downto 0);
	signal RoundKey								: STD_LOGIC_VECTOR(63 downto 0);
	signal CiphertextRegIn						: STD_LOGIC_VECTOR(63 downto 0);
	
	signal K0										: STD_LOGIC_VECTOR(63 downto 0);
	signal K1										: STD_LOGIC_VECTOR(63 downto 0);
	
	signal FSM										: STD_LOGIC_VECTOR(5  downto 0);
	signal FSMUpdate								: STD_LOGIC_VECTOR(5  downto 0);
	signal FSMSelected							: STD_LOGIC_VECTOR(5  downto 0);
	signal AddKey									: STD_LOGIC_VECTOR(0  downto 0);
	signal SelKey									: STD_LOGIC_VECTOR(0  downto 0);
	signal done_internal							: STD_LOGIC_VECTOR(0  downto 0);

	------

	signal Red_Plaintext							: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);
	signal Red_StateRegOutput					: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);
	signal Red_StateRegInput					: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);
	signal Red_AddRoundKeyOutput				: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);
	signal Red_AddKeyMUXOutput					: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);
	signal Red_AddConstInput					: STD_LOGIC_VECTOR(8*Red_size-1  downto 0);
	signal Red_AddConstOutput					: STD_LOGIC_VECTOR(8*Red_size-1  downto 0);	
	signal Red_AddConstMUXOutput					: STD_LOGIC_VECTOR(8*Red_size-1  downto 0);
	signal Red_ShiftRowsInput					: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);
	signal Red_Feedback							: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);
	signal Red_RoundKey							: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);

	signal Red_K0									: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);
	signal Red_K1									: STD_LOGIC_VECTOR(16*Red_size-1 downto 0);

	signal Error									: STD_LOGIC_VECTOR(Red_size-1   downto 0);
	signal ErrorFree								: STD_LOGIC_VECTOR(Error_size-1 downto 0);
	signal ErrorFreeUpdate						: STD_LOGIC_VECTOR(Error_size-1 downto 0);

	signal Red_AddKey								: STD_LOGIC_VECTOR(Red_size-1 downto 0);
	signal Red_SelKey								: STD_LOGIC_VECTOR(Red_size-1 downto 0);
	signal Red_done								: STD_LOGIC_VECTOR(Red_size-1 downto 0);

	signal SignaltoCheck							: STD_LOGIC_VECTOR(ToCheckCount*4-1 downto 0);
	signal Red_SignaltoCheck					: STD_LOGIC_VECTOR(ToCheckCount*Red_size-1 downto 0);
	signal Red_final								: STD_LOGIC_VECTOR(ToCheckCount*Red_size-1 downto 0);

	signal Red_FSM									: STD_LOGIC_VECTOR(2*Red_size-1 downto 0);
	signal Red_FSMUpdate							: STD_LOGIC_VECTOR(2*Red_size-1 downto 0);
	signal Red_FSMSelected						: STD_LOGIC_VECTOR(2*Red_size-1 downto 0);
	signal Red_FSMStart						   : STD_LOGIC_VECTOR(2*Red_size-1 downto 0);
	
begin

	PlaintextMUX: ENTITY work.MUX
	GENERIC Map ( size => 64)
	PORT Map ( 
		sel	=> rst,
		D0   	=> Feedback,
		D1 	=> Plaintext,
		Q 		=> StateRegInput);

	StateReg: ENTITY work.reg
	GENERIC Map ( size => 64)
	PORT Map ( 
		clk	=> clk,
		D 		=> StateRegInput,
		Q 		=> StateRegOutput);

	AddKeyXOR: ENTITY work.XOR_2n
	GENERIC Map ( size => 4, count => 16)
	PORT Map ( StateRegOutput, RoundKey, AddRoundKeyOutput);

	AddKeyMUX: ENTITY work.MUX
	GENERIC Map ( size => 64)
	PORT Map ( 
		sel	=> AddKey(0),
		D0   	=> StateRegOutput,
		D1 	=> AddRoundKeyOutput,
		Q 		=> AddKeyMUXOutput);

	AddConstInput  <= AddKeyMUXOutput(63 downto 56) & AddKeyMUXOutput(47 downto 40) & AddKeyMUXOutput(31 downto 24) & AddKeyMUXOutput(15 downto 8);
	AddConstInput2 <= '0' & FSM(5 downto 3) & '0' & FSM(2 downto 0);
	
	AddConstXOR: ENTITY work.AddConst
	GENERIC Map ( 4, Identity, x"0")
	PORT Map ( AddConstInput, AddConstInput2, AddConstOutput);

	AddConstMUX: ENTITY work.MUX
	GENERIC Map ( size => 32)
	PORT Map ( 
		sel	=> done_internal(0),
		D0   	=> AddConstOutput,
		D1 	=> AddConstInput,
		Q 		=> AddConstMUXOutput);

	ShiftRowsInput <= AddConstMUXOutput(31 downto 24) & AddKeyMUXOutput(55 downto 48) &
	                  AddConstMUXOutput(23 downto 16) & AddKeyMUXOutput(39 downto 32) &
						   AddConstMUXOutput(15 downto 8)  & AddKeyMUXOutput(23 downto 16) &
						   AddConstMUXOutput(7  downto 0)  & AddKeyMUXOutput(7  downto 0);

	ShiftRowsInst: ENTITY work.ShiftRows
	GENERIC Map ( size => 4)
	PORT Map (
		state		=> ShiftRowsInput,
		result	=> ShiftRowsOutput);
		
	MCInst: ENTITY work.SB_MC
	GENERIC Map ( SboxTable, 4, Identity, x"0")
	PORT Map (
		state		=> ShiftRowsOutput,
		result	=> Feedback);

	-----------------------------------------------	
	
	Red_PlaintextInst: ENTITY work.FMulti
	GENERIC Map ( size => Red_size, count => 16, Table => LFTable)
	PORT Map (
		input		=> Plaintext,
		output	=> Red_Plaintext);
		
	Red_PlaintextMUX: ENTITY work.MUX
	GENERIC Map ( size => 16*Red_size)
	PORT Map ( 
		sel	=> rst,
		D0		=> Red_Feedback,
		D1		=> Red_Plaintext,
		Q		=> Red_StateRegInput);

	Red_StateReg: ENTITY work.reg
	GENERIC Map ( size => Red_size*16)
	PORT Map ( 
		clk	=> clk,
		D 		=> Red_StateRegInput,
		Q 		=> Red_StateRegOutput);
		
	RedAddKeyXOR: ENTITY work.XOR_2n
	GENERIC Map ( size => Red_size, count => 16)
	PORT Map ( Red_StateRegOutput, Red_RoundKey, Red_AddRoundKeyOutput, LFC(Red_size-1 downto 0));

	RedAddKeyMUX: ENTITY work.MUX2to1_Redn
	GENERIC Map ( 
		size1   => Red_size, 
		size2   => 16*Red_size,
		LFTable => LFTable)
	PORT Map ( 
		sel	=> Red_AddKey,
		D0   	=> Red_StateRegOutput,
		D1 	=> Red_AddRoundKeyOutput,
		Q 		=> Red_AddKeyMUXOutput);
		
	Red_AddConstInput <= Red_AddKeyMUXOutput(Red_size*16-1 downto Red_size*14) & 
								Red_AddKeyMUXOutput(Red_size*12-1 downto Red_size*10) & 
								Red_AddKeyMUXOutput(Red_size*8-1  downto Red_size*6) & 
								Red_AddKeyMUXOutput(Red_size*4-1  downto Red_size*2);

	Red_AddConstXOR: ENTITY work.AddConst
	GENERIC Map (Red_size, LFTable, LFC)
	PORT Map ( Red_AddConstInput, Red_FSM, Red_AddConstOutput);

	RedAddConstMUX: ENTITY work.MUX2to1_Redn
	GENERIC Map ( 
		size1   => Red_size, 
		size2   => 8*Red_size,
		LFTable => LFTable)
	PORT Map ( 
		sel	=> Red_done,
		D0   	=> Red_AddConstOutput,
		D1 	=> Red_AddConstInput,
		Q 		=> Red_AddConstMUXOutput);

	Red_ShiftRowsInput <= Red_AddConstMUXOutput(Red_size*8-1 downto Red_size*6) & Red_AddKeyMUXOutput(Red_size*14-1 downto Red_size*12) &
							    Red_AddConstMUXOutput(Red_size*6-1 downto Red_size*4) & Red_AddKeyMUXOutput(Red_size*10-1 downto Red_size*8) &
							    Red_AddConstMUXOutput(Red_size*4-1 downto Red_size*2) & Red_AddKeyMUXOutput(Red_size*6-1  downto Red_size*4) &
							    Red_AddConstMUXOutput(Red_size*2-1 downto 0)          & Red_AddKeyMUXOutput(Red_size*2-1  downto 0);

	----	
		
	Red_MCInst: ENTITY work.SB_MC
	GENERIC Map ( SboxTable, Red_size, LFTable, LFC)
	PORT Map (
		state		=> ShiftRowsOutput,
		result	=> Red_Feedback);
		
	--===================================================

	K0		<= Key(127 downto 64);
	K1		<= Key( 63 downto  0);

	KeyMUX: ENTITY work.MUX
	GENERIC Map ( size => 64)
	PORT Map ( 
		sel	=> SelKey(0),
		D0   	=> K0,
		D1 	=> K1,
		Q 		=> RoundKey);	
	
	--------------------------
	
	Red_K0Inst: ENTITY work.FMulti
	GENERIC Map ( size => Red_size, count => 16, Table => LFTable)
	PORT Map (
		input		=> K0,
		output	=> Red_K0);
		
	Red_K1Inst: ENTITY work.FMulti
	GENERIC Map ( size => Red_size, count => 16, Table => LFTable)
	PORT Map (
		input		=> K1,
		output	=> Red_K1);
	
	Red_KeyMUX: ENTITY work.MUX2to1_Redn
	GENERIC Map ( 
		size1   => Red_size,
		size2   => 16*Red_size,
		LFTable => LFTable)
	PORT Map (
		sel	=> Red_SelKey,
		D0		=> Red_K0,
		D1		=> Red_K1,
		Q		=> Red_RoundKey);	
		
	-----------------------------------------------
	
	GENMV0:
	IF MultiVariate = 0 GENERATE
		SignaltoCheck <= "000" & done_internal & "000" & AddKey & "000" & SelKey & '0' & FSM(5 downto 3) & '0' & FSM(2 downto 0) & ShiftRowsInput;
		Red_final     <= Red_done & Red_AddKey & Red_SelKey & Red_FSM & Red_ShiftRowsInput;
	END GENERATE;
	
	GENMV1:
	IF MultiVariate = 1 GENERATE
		SignaltoCheck <= "000" & done_internal & "000" & AddKey & "000" & SelKey & '0' & FSM(5 downto 3) & '0' & FSM(2 downto 0) & ShiftRowsInput &
		                 '0' & FSMSelected(5 downto 3) & '0' & FSMSelected(2 downto 0) & StateRegInput;
		Red_final     <= Red_done & Red_AddKey & Red_SelKey & Red_FSM & Red_ShiftRowsInput &
				           Red_FSMSelected & Red_StateRegInput;
	END GENERATE;

	--------
	
	Red_ToCheckInst: ENTITY work.FMulti
		GENERIC Map ( size  => Red_size, count => ToCheckCount, Table => LFTable)
		PORT Map (
			input		=> SignaltoCheck,
			output	=> Red_SignaltoCheck);
		
	Check1: ENTITY work.Checkn
	GENERIC Map ( count => ToCheckCount, sizecount => 1, size  => Red_size)
	PORT Map ( 
		in1		=> Red_final,
		in2    	=> Red_SignaltoCheck,
		result 	=> Error);
		
	-------------------------------------
	
	GEN1 :
	FOR i IN 0 TO Error_size-1 GENERATE
		ANDInst: ENTITY work.ANDn
		Generic Map (size1 => Red_size, size2 => Error_size)
		Port Map (Error, ErrorFree, ErrorFreeUpdate(i));
	END GENERATE;

	ErrorDetectionReg: PROCESS(clk, rst, ErrorFreeUpdate)
	BEGIN
		IF RISING_EDGE(clk) THEN
			IF (rst = '1') THEN
				ErrorFree	<= (others => '1');
			ELSE
				ErrorFree 	<= ErrorFreeUpdate;
			END IF;
		END IF;
	END PROCESS;		
		
	--------------
	
	OutputMUX: ENTITY work.MUX2to1_Redn_forcheck
	GENERIC Map ( 
		size1   => Error_size,
		size2	  => 64)
	PORT Map (
		sel	=> ErrorFreeUpdate,
		D0		=> (others => '0'),
		D1		=> ShiftRowsInput,
		Q		=> CiphertextRegIn);
				
	CiphertextReg: ENTITY work.regER
	GENERIC Map ( size => 64)
	PORT Map ( 
		clk	=> clk,
		rst	=> rst,
		EN		=> done_internal(0),
		D 		=> CiphertextRegIn,
		Q 		=> Ciphertext);

	-------------------------------------
	
	FSMMUX: ENTITY work.MUX
	GENERIC Map ( size => 6)
	PORT Map ( 
		sel	=> rst,
		D0   	=> FSMUpdate,
		D1 	=> "000001",
		Q 		=> FSMSelected);
		
	FSMReg: ENTITY work.reg
	GENERIC Map ( size => 6)
	PORT Map ( 
		clk	=> clk,
		D 		=> FSMSelected,
		Q 		=> FSM);
		
	FSMUpdateInst: ENTITY work.StateUpdate
	GENERIC Map ( 3, Identity )
	PORT Map (FSM, FSMUpdate);
	
	FSMSignalsInst: ENTITY work.FSMSignals
	GENERIC Map ( 1, Identity )
	PORT Map (FSM, AddKey, SelKey, done_internal);

	----------------
	
	Red_FSMStart <= LFTable(60+Red_size-1 downto 60) & LFTable(56+Red_size-1 downto 56); -- LF( 0000) & LF(0001)
	
	Red_FSMMUX: ENTITY work.MUX
	GENERIC Map ( size => 2*Red_size)
	PORT Map ( 
		sel	=> rst,
		D0		=> Red_FSMUpdate,
		D1		=> Red_FSMStart,
		Q		=> Red_FSMSelected);		
		
	Red_FSMReg: ENTITY work.reg
	GENERIC Map ( size => 2*Red_size)
	PORT Map ( 
		clk	=> clk,
		D 		=> Red_FSMSelected,
		Q 		=> Red_FSM);
	
	Red_FSMUpdateInst: ENTITY work.StateUpdate
	GENERIC Map ( Red_size, LFTable )
	PORT Map (FSM, Red_FSMUpdate);
	
	Red_FSMSignalsInst: ENTITY work.FSMSignals
	GENERIC Map ( Red_size, LFTable )
	PORT Map (FSM, Red_AddKey, Red_SelKey, Red_done);

	done		<= done_internal(0);	

end Behavioral;

