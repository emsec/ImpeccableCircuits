----------------------------------------------------------------------------------
-- COMPANY:		Ruhr University Bochum, Embedded Security
-- AUTHOR:		https://eprint.iacr.org/2018/203
----------------------------------------------------------------------------------
-- Copyright (c) 2019, Anita Aghaie, Amir Moradi
-- All rights reserved.

-- BSD-3-Clause License
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--     * Redistributions of source code must retain the above copyright
--       notice, this list of conditions and the following disclaimer.
--     * Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
--     * Neither the name of the copyright holder, their organization nor the
--       names of its contributors may be used to endorse or promote products
--       derived from this software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;
use work.functions.all;

entity FSMSignals is
    Port ( FSM   		: in   STD_LOGIC_VECTOR (4 downto 0);
           last  		: out  STD_LOGIC;
			  done  		: out  STD_LOGIC;
			  sel_K0_1	: out  STD_LOGIC;
			  sel_K_WK	: out  STD_LOGIC);
end FSMSignals;

architecture Behavioral of FSMSignals is
begin

	lastInst: ENTITY work.LookUp
	GENERIC Map (size => 5, Table => MakeSignallastTable)
	PORT Map (FSM, last);

	doneInst: ENTITY work.LookUp
	GENERIC Map (size => 5, Table => MakeSignaldoneTable)
	PORT Map (FSM, done);

	sel_K0_1Inst: ENTITY work.LookUp
	GENERIC Map (size => 5, Table => MakeSignalsel_K0_1Table)
	PORT Map (FSM, sel_K0_1);

	sel_K_WKInst: ENTITY work.LookUp
	GENERIC Map (size => 5, Table => MakeSignalsel_K_WKTable)
	PORT Map (FSM, sel_K_WK);

end Behavioral;

