----------------------------------------------------------------------------------
-- COMPANY:		Ruhr University Bochum, Embedded Security
-- AUTHOR:		https://eprint.iacr.org/2018/203
----------------------------------------------------------------------------------
-- Copyright (c) 2019, Amir Moradi, Aein Rezaei Shahmirzadi
-- All rights reserved.

-- BSD-3-Clause License
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--     * Redistributions of source code must retain the above copyright
--       notice, this list of conditions and the following disclaimer.
--     * Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
--     * Neither the name of the copyright holder, their organization nor the
--       names of its contributors may be used to endorse or promote products
--       derived from this software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity RconFSM is
    Port ( clk : in  STD_LOGIC;
			  rst : in  STD_LOGIC;
           InitialRound : out  STD_LOGIC;
           FinalRound : out  STD_LOGIC;
			  done : out  STD_LOGIC;
           rcon : out  STD_LOGIC_VECTOR (7 downto 0));
end RconFSM;

architecture Behavioral of RconFSM is

	signal RegIn, RegOut, Xor2In, conditionalXOR : STD_LOGIC_VECTOR (7 DOWNTO 0);

begin

	StateRegR: ENTITY work.regR 
	GENERIC Map ( size => 8)
	PORT MAP(
		clk => clk,
		rst => rst,
		D => RegIn,
		Q => RegOut);
	
	Xor2In 			<= RegOut(6 downto 0) & "0";
	conditionalXOR <= "000" & RegOut(7) & RegOut(7) & "0" & RegOut(7) & RegOut(7);
	
	rcon_XOR2: ENTITY work.XOR_2n
	GENERIC Map ( size => 8, count => 1)
	PORT Map ( Xor2In, conditionalXOR, RegIn);

	rcon <= RegOut;
	
	FSM_Gen: PROCESS(RegOut)
	BEGIN
		
		IF (RegOut = x"01") THEN
			InitialRound	<= '1';
		ELSE 
			InitialRound	<= '0';
		END IF;
		
		IF (RegOut = x"6c") THEN
			FinalRound	<= '1';
		ELSE 
			FinalRound	<= '0';
		END IF;
		
		IF (RegOut = x"d8") THEN
			done	<= '1';
		ELSE 
			done	<= '0';
		END IF;
	
	END PROCESS;
	
end Behavioral;

