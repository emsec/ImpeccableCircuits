----------------------------------------------------------------------------------
-- COMPANY:		Ruhr University Bochum, Embedded Security
-- AUTHOR:		https://eprint.iacr.org/2018/203
----------------------------------------------------------------------------------
-- Copyright (c) 2019, Anita Aghaie, Amir Moradi
-- All rights reserved.

-- BSD-3-Clause License
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--     * Redistributions of source code must retain the above copyright
--       notice, this list of conditions and the following disclaimer.
--     * Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
--     * Neither the name of the copyright holder, their organization nor the
--       names of its contributors may be used to endorse or promote products
--       derived from this software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY RoundConstant_MUX IS
	PORT ( Round : IN  STD_LOGIC_VECTOR (3 DOWNTO 0);
			 RoundConstant : OUT  STD_LOGIC_VECTOR (63 DOWNTO 0));
END RoundConstant_MUX;

ARCHITECTURE behavioral OF RoundConstant_MUX IS

	signal RCLSB	: std_logic_vector(15 downto 0);

BEGIN

	RCInst: ENTITY work.RoundConstant
	PORT Map ( 
		Round  => Round,
		RCLSB  => RCLSB);

	RoundConstant	<= "000" & RCLSB(15) & "000" & RCLSB(14) & "000" & RCLSB(13) & "000" & RCLSB(12) & 
	                  "000" & RCLSB(11) & "000" & RCLSB(10) & "000" & RCLSB(9) & "000" & RCLSB(8) & 
							"000" & RCLSB(7) & "000" & RCLSB(6) & "000" & RCLSB(5) & "000" & RCLSB(4) & 
							"000" & RCLSB(3) & "000" & RCLSB(2) & "000" & RCLSB(1) & "000" & RCLSB(0);

END behavioral;

