----------------------------------------------------------------------------------
-- COMPANY:		Ruhr University Bochum, Embedded Security
-- AUTHOR:		https://doi.org/10.13154/tosc.v2019.i1.5-45 
----------------------------------------------------------------------------------
-- Copyright (c) 2019, Amir Moradi 
-- All rights reserved.

-- BSD-3-Clause License
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--     * Redistributions of source code must retain the above copyright
--       notice, this list of conditions and the following disclaimer.
--     * Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
--     * Neither the name of the copyright holder, their organization nor the
--       names of its contributors may be used to endorse or promote products
--       derived from this software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity selectsUpdateBit is
	Generic (withDec			: integer;
				BitNumber   	: integer);
	Port ( selects   			: in  STD_LOGIC_VECTOR (1 downto 0);
			 FSM3					: in  STD_LOGIC;
			 EncDec	  			: in  STD_LOGIC;
          selectsNextBit	: out STD_LOGIC);
end selectsUpdateBit;

architecture Behavioral of selectsUpdateBit is
begin

	GEN0: IF BitNumber=0 GENERATE
		selectsNextBit		<= selects(0) XOR FSM3;
	END GENERATE;	
	
	GEN1: IF BitNumber=1 GENERATE
		GenwithoutDecselects: IF withDec = 0 GENERATE
			selectsNextBit		<= selects(1) XOR (FSM3 AND selects(0));
		END GENERATE;
		
		GenwithDecselects: IF withDec /= 0 GENERATE
			selectsNextBit		<= selects(1) XOR (FSM3 AND (selects(0) XOR EncDec));
		END GENERATE;
	END GENERATE;	

end Behavioral;


