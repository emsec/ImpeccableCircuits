----------------------------------------------------------------------------------
-- COMPANY:		Ruhr University Bochum, Embedded Security
-- AUTHOR:		https://eprint.iacr.org/2018/203
----------------------------------------------------------------------------------
-- Copyright (c) 2019, Anita Aghaie, Amir Moradi, Aein Rezaei Shahmirzadi
-- All rights reserved.

-- BSD-3-Clause License
-- Redistribution and use in source and binary forms, with or without
-- modification, are permitted provided that the following conditions are met:
--     * Redistributions of source code must retain the above copyright
--       notice, this list of conditions and the following disclaimer.
--     * Redistributions in binary form must reproduce the above copyright
--       notice, this list of conditions and the following disclaimer in the
--       documentation and/or other materials provided with the distribution.
--     * Neither the name of the copyright holder, their organization nor the
--       names of its contributors may be used to endorse or promote products
--       derived from this software without specific prior written permission.
-- 
-- THIS SOFTWARE IS PROVIDED BY THE COPYRIGHT HOLDERS AND CONTRIBUTORS "AS IS" AND
-- ANY EXPRESS OR IMPLIED WARRANTIES, INCLUDING, BUT NOT LIMITED TO, THE IMPLIED
-- WARRANTIES OF MERCHANTABILITY AND FITNESS FOR A PARTICULAR PURPOSE ARE
-- DISCLAIMED. IN NO EVENT SHALL THE COPYRIGHT HOLDER OR CONTRIBUTERS BE LIABLE FOR ANY
-- DIRECT, INDIRECT, INCIDENTAL, SPECIAL, EXEMPLARY, OR CONSEQUENTIAL DAMAGES
-- (INCLUDING, BUT NOT LIMITED TO, PROCUREMENT OF SUBSTITUTE GOODS OR SERVICES;
-- LOSS OF USE, DATA, OR PROFITS; OR BUSINESS INTERRUPTION) HOWEVER CAUSED AND
-- ON ANY THEORY OF LIABILITY, WHETHER IN CONTRACT, STRICT LIABILITY, OR TORT
-- (INCLUDING NEGLIGENCE OR OTHERWISE) ARISING IN ANY WAY OUT OF THE USE OF THIS
-- SOFTWARE, EVEN IF ADVISED OF THE POSSIBILITY OF SUCH DAMAGE.

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

ENTITY RedMC IS
	generic(Red_size : positive;
			  Table : STD_LOGIC_VECTOR (2047 DOWNTO 0));
	PORT ( data_in  : IN  STD_LOGIC_VECTOR (127 DOWNTO 0);
			 Red_in	 : IN  STD_LOGIC_VECTOR (Red_size*16-1 DOWNTO 0);		
			 data_out : OUT STD_LOGIC_VECTOR (Red_size*16-1 DOWNTO 0));		
END RedMC;

ARCHITECTURE behavioral OF RedMC IS	

BEGIN

	GEN :
	FOR i IN 0 TO 3 GENERATE
		Inst_RedMixOneColumn: ENTITY work.RedMixOneColumn
		GENERIC Map ( Red_size => Red_size, Table => Table)
		PORT MAP(
			data_in  => data_in((i+1)*32-1 downto i*32),
			Red_in   => Red_in  ((i+1)*Red_size*4-1 downto i*Red_size*4),
			data_out => data_out((i+1)*Red_size*4-1 downto i*Red_size*4));
	END GENERATE;

END behavioral;

